`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Electronics Corporation of India Limited
// Engineer: Rishav Ambasta
// 
// Create Date:    19:33:17 07/02/2014 
// Design Name: 
// Module Name:    Rx 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Rx(
    );


endmodule
